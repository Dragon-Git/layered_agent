package up_agt_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "up_item.sv"
    `include "up_drv.sv"
    `include "up_sqr.sv"
    `include "up_agt.sv"
    // `include "up_reg_adapter.sv"

endpackage: up_agt_pkg