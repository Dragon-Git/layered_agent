package typical_env_pkg;
    import uvm_pkg::*;  
    `include "uvm_macros.svh"

    import up_agt_pkg::*;
    import regmap_pkg::*;

    `include "reg_item.sv"
    `include "reg_adapter.sv"
    `include "reg_adapter_seq.sv"
    `include "base_env.sv"
    `include "base_test.sv"

endpackage: typical_env_pkg
